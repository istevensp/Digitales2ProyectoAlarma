veinte5_inst : veinte5 PORT MAP (
		result	 => result_sig
	);
