diez4_inst : diez4 PORT MAP (
		result	 => result_sig
	);
