num_k_inst : num_k PORT MAP (
		result	 => result_sig
	);
