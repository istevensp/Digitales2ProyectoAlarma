nueve4_inst : nueve4 PORT MAP (
		result	 => result_sig
	);
