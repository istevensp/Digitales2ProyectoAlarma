num_i_inst : num_i PORT MAP (
		result	 => result_sig
	);
