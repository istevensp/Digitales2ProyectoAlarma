seis4_inst : seis4 PORT MAP (
		result	 => result_sig
	);
