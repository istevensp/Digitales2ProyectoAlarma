tres4_inst : tres4 PORT MAP (
		result	 => result_sig
	);
