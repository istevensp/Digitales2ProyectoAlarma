siete4_inst : siete4 PORT MAP (
		result	 => result_sig
	);
