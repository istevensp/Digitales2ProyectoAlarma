ocho4_inst : ocho4 PORT MAP (
		result	 => result_sig
	);
