uno4_inst : uno4 PORT MAP (
		result	 => result_sig
	);
