cinco4_inst : cinco4 PORT MAP (
		result	 => result_sig
	);
