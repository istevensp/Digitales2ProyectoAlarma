num_j_inst : num_j PORT MAP (
		result	 => result_sig
	);
